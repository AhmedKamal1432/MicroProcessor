library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


Entity Control_Store is
  port(
    Rst,clk : in std_logic;
    Add:in std_logic_vector(7 downto 0);
    Control_Word:out std_logic_vector(31 downto 0));  
end Control_Store;

architecture Control_Store of Control_Store is
  type ram_type is array(0 to 1024) of std_logic_vector(31 downto 0);

  signal rom : ram_type := ( 
    000 =>  "00000001000101101000001011100000", 
    001 =>  "00000010001100100000000000000000", 
    002 =>  "00000011001001000000000000000000", 
    003 =>  "00000000000000000000000000000001", 
    4   =>  "00000000000000000000000110000000",
    16  =>  "10111100100001100000001001011000",
    17  =>  "10111100100001100000001000011000",
    18  =>  "10111100100001100000010000111000",
    20  =>  "00011101000000000000000000000000",
    21  =>  "10111100100001100000101000011000",
    22  =>  "10111100100001100000110000011000",
    23  =>  "00011000000001100000000000000000",
    24  =>  "00011001001100011000000000000000",
    25  =>  "00011010100000000010000000000000",
    26  =>  "00000000101000000000010000110000",
    28  =>  "00000000100000000000100000010000",
    29  =>  "00011110000001100000000000000000",
    30  =>  "00011111001100011000000000000000",
    31  =>  "00100000100000000010000000000000",
    32  =>  "00100001000001100000111000000000",
    33  =>  "00100010001100000010000000000000",
    34  =>  "10111100101001100000100000011000",
    65  =>  "10000001010000000100000000000010",
    73  =>  "01001010010000001000000010000000",
    74  =>  "01111001000000000000000000000000",
    81  =>  "01010010010001101000001011100000",
    82  =>  "01111000001110000000000000000100",
    97  =>  "01100010010000000010000000000000",
    98  =>  "01100011000001100000011000000000",
    99  =>  "01100100001110001000000010000000",
    100 =>  "01111000000000000000000000000100",
    113 =>  "01110010000101101000001011100000",
    114 =>  "01110011001100100000000000000000",
    115 =>  "01110100001000000010000000000000",
    116 =>  "01110101010001100000001000000000",
    117 =>  "01110110001100001000000010000000",
    118 =>  "01111000000000000000000000000100",
    120 =>  "00000110001000001000000010000000",
    6   =>  "01111001000000000000000000000000",
    121 =>  "10000001001000000100000000000010",
    129 =>  "00010000010100000010000000001010",
    137 =>  "10001010010100001000000010000000",
    138 =>  "10111001000000000000000000000000",
    145 =>  "10010010010101101000001011100000",
    146 =>  "10111000001110100000000000000110",
    161 =>  "10100010010100000010000000000000",
    162 =>  "10100011000001100000011000000000",
    163 =>  "10100100001110101000000010000000",
    164 =>  "10111000000000000000000000000110",
    177 =>  "10110010000101101000001011100000",
    178 =>  "10110011001100100000000000000000",
    179 =>  "10110100001000000010000000000000",
    180 =>  "10110101010101100000001000000000",
    181 =>  "10110110001100001000000010000000",
    182 =>  "10111000000000000000000000000110",
    184 =>  "00000111001000001000000010000000",
    7   =>  "10111001000000000000000000000000",
    185 =>  "00010000001000000010000000001010",
    188 =>  "00000000001100010000000100000000",
    189 =>  "00000000001110100000000000000000",
  others => "00000000000000000000000000000000"   
  );

begin
 process(clk,Rst) is
    Begin
    if Rst='1' then
       Control_Word<=(others=>'0');
    elsif falling_edge(clk) and  Rst='0' then  
      Control_Word <= rom(to_integer(unsigned(Add)));

    end if;
  end process;
end Control_Store;
