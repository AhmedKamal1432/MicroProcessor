library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


Entity Control_Store is
  port(
    Rst,clk : in std_logic;
    Add:in std_logic_vector(7 downto 0);
    Control_Word:out std_logic_vector(31 downto 0));  
end Control_Store;

architecture Control_Store of Control_Store is
  type ram_type is array(0 to 1024) of std_logic_vector(31 downto 0);

  signal rom : ram_type := ( 
  0   => "00000001000101101000001011100000", 
  1   => "00000010001100100000000000000000", 
  2   => "00000011001001000000000000000000", 
  3   => "00000000000000000000000000000001", 
4	=>	"00000000000000000000000110000000",
16	=>	"10111100100001100000001001011000",
17	=>	"10111100100001100000001000011000",
18	=>	"10111100100001100000010000111000",
20	=>	"00011101000000000000000000000000",
21	=>	"10111100100001100000101000011000",
22	=>	"10111100100001100000110000011000",
23	=>	"00011000000001100000000000000000",
24	=>	"00011001001100011000000000000000",
25	=>	"00011010100000000010000000000000",
26	=>	"00000000101000000000010000110000",
28	=>	"00000000100000000000100000010000",
29	=>	"00011110000001100000000000000000",
30	=>	"00011111001100011000000000000000",
31	=>	"00100000100000000010000000000000",
32	=>	"00100001000001100000111000000000",
33	=>	"00100010001100000010000000000000",
34	=>	"10111100101001100000100000011000",
65	=>	"10000001010000000100000000000010",
73	=>	"01001010010000001000000010000000",
74	=>	"01111001000000000000000000000000",
81	=>	"01010010010001101000001011100000",
82	=>	"01111000001110000000000000000100",
97	=>	"01100010010000000010000000000000",
98	=>	"01100011000001100000011000000000",
99	=>	"01100100001110001000000010000000",
100	=>	"01111000000000000000000000000100",
113	=>	"01110010000101101000001011100000",
114	=>	"01110011001100100000000000000000",
115	=>	"01110100001000000010000000000000",
116	=>	"01110101010001100000001000000000",
117	=>	"01110110001100001000000010000000",
118	=>	"01111000000000000000000000000100",
120	=>	"10000010001000001000000010000000",
130	=>	"01111001000000000000000000000000",
121	=>	"10000001001000000100000000000010",
129	=>	"00000000010100000010000000001010",
137	=>	"10001010010100001000000010000000",
138	=>	"10111001000000000000000000000000",
145	=>	"10010010010101101000001011100000",
146	=>	"10111000001110100000000000000110",
161	=>	"10100010010100000010000000000000",
162	=>	"10100011000001100000011000000000",
163	=>	"10100100001110101000000010000000",
164	=>	"10111000000000000000000000000110",
177	=>	"10110010000101101000001011100000",
178	=>	"10110011001100100000000000000000",
179	=>	"10110100001000000010000000000000",
180	=>	"10110101010101100000001000000000",
181	=>	"10110110001100001000000010000000",
182	=>	"10111000000000000000000000000110",
184	=>	"10000011001000001000000010000000",
131	=>	"10111001000000000000000000000000",
185	=>	"00000000001000000010000000001010",
188	=>	"00000000001100010000000100000000",
189	=>	"00000000001110100000000000000000",
48	=>	"00110100000000000000000000001100",
51	=>	"00000110000000000000000000001100",
52	=>	"10111100000001100000000000111000",
53	=>	"00110110000001100000000000000000",
54	=>	"00000000001100100000000000000000",
6	=>	"10111100000001100000011000011000",
7	=>	"10111100000001100000011000111000",
55	=>	"10111100000001100000111000011000",
56	=>	"10111100000001100001000000011000",
57	=>	"10111100000001100001001000011000",
58	=>	"10111100000001100001010000011000",
59	=>	"10111100000001100001011000011000",
60	=>	"10111100000001100001100000011000",
61	=>	"10111100000001100001101000011000",
62	=>	"10111100000001100001110000011000",
63	=>	"10111100000001100001111000011000",
140	=>	"10001101000100000010000000000000",
141	=>	"10001110101101100000001000000000",
142	=>	"00000000001100100000000000000000",
8	=>	"00001001000001100000000000000000",
9	=>	"00001010001100011000000000000000",
10	=>	"00001011110000000010000000000000",
11	=>	"00001100000001100000011000000000",
12	=>	"00001101001111001000000000000000",
13	=>	"00001110010000010000000100000000",
14	=>	"00001111000110000000000000000000",
15	=>	"00000000101000100000000000000000",
75	=>	"01001100010000100000000000000000",
76	=>	"01001101110000001010000010000000",
77	=>	"01001110000001100000000000100000",
78	=>	"01001111001010000000000000000000",
79	=>	"00000000001111000000000000000000",
 others => "00000000000000000000000000000000"   
  );

begin
 process(clk,Rst) is
    Begin
    if Rst='1' then
       Control_Word<=(others=>'0');
    elsif falling_edge(clk) and  Rst='0' then  
      Control_Word <= rom(to_integer(unsigned(Add)));

    end if;
  end process;
end Control_Store;
